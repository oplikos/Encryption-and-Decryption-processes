// Code your design here
`include "Definitions.sv"
`include "InstFetch.sv"
`include "ALU.sv"
`include "Ctrl.sv"
`include "DataMem.sv"
`include "top_level.sv"
`include "Immediate_LUT.sv"
`include "InstROM.sv"
`include "RegFile.sv"
`include "Mux.sv"