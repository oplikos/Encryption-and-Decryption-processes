// Code your testbench here
// or browse Examples
//`include "program1_tb1.sv"
`include "program2.sv"
//`include "program3.sv"